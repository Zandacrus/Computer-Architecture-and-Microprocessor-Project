/*
	Arkanil
*/